/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: comparator 
-----------------------------------------------------------*/
`timescale 1 ns/1 ns
module comparator(
 category,
 overweight,
 normal,
 underweight);
  input [7:0] category;
  output overweight;
  output normal;
  output underweight;
 // write your code here, please.
endmodule